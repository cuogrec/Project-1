library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity sine_lut is
    port(
        fsclk  : in  std_logic;
        rst    : in  std_logic;
        data_o : out std_logic_vector(11 downto 0)
    );
end entity;

architecture rtl of sine_lut is
    type rom_t is array(0 to 63) of std_logic_vector(11 downto 0);
    constant ROM : rom_t := (
        0  => "100000000000",
        1  => "100011001001",
        2  => "100110001111",
        3  => "101001010010",
        4  => "101100001111",
        5  => "101111000101",
        6  => "110001110001",
        7  => "110100010011",
        8  => "110110101000",
        9  => "111000101111",
        10 => "111010100111",
        11 => "111100001110",
        12 => "111101100100",
        13 => "111110100111",
        14 => "111111011000",
        15 => "111111110110",
        16 => "111111111111",
        17 => "111111110110",
        18 => "111111011000",
        19 => "111110100111",
        20 => "111101100100",
        21 => "111100001110",
        22 => "111010100111",
        23 => "111000101111",
        24 => "110110101000",
        25 => "110100010011",
        26 => "110001110001",
        27 => "101111000101",
        28 => "101100001111",
        29 => "101001010010",
        30 => "100110001111",
        31 => "100011001001",
        32 => "100000000000",
        33 => "011100110111",
        34 => "011001110001",
        35 => "010110101110",
        36 => "010011110001",
        37 => "010000111011",
        38 => "001110001111",
        39 => "001011101101",
        40 => "001001010000",
        41 => "000111001001",
        42 => "000101010001",
        43 => "000011101010",
        44 => "000010010100",
        45 => "000001010001",
        46 => "000000100000",
        47 => "000000000010",
        48 => "000000000000",
        49 => "000000000010",
        50 => "000000100000",
        51 => "000001010001",
        52 => "000010010100",
        53 => "000011101010",
        54 => "000101010001",
        55 => "000111001001",
        56 => "001001010000",
        57 => "001011101101",
        58 => "001110001111",
        59 => "010000111011",
        60 => "010011110001",
        61 => "010110101110",
        62 => "011001110001",
        63 => "011100110111"
    );

    signal addr : unsigned(5 downto 0) := (others=>'0');
begin
    process(fsclk)
    begin
        if rising_edge(fsclk) then
            if rst='1' then
                addr <= (others=>'0');
            else
                addr <= addr + 1;
            end if;
        end if;
    end process;

    data_o <= ROM(to_integer(addr));
end architecture;
